interface intf();
  logic [3:0]a,b,s;
  logic cy;
endinterface