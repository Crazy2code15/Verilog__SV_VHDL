interface intf();
  logic a,b,cin,s,cy;
endinterface